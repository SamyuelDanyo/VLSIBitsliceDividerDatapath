magic
tech c35b4
timestamp 1543772130
<< pimplant >>
rect 0 334 252 727
<< nimplant >>
rect 0 31 252 281
<< nwell >>
rect 0 334 252 752
<< polysilicon >>
rect 188 710 195 718
rect 216 710 223 718
rect 46 692 53 701
rect 73 692 80 701
rect 126 692 133 701
rect 46 624 53 636
rect 73 624 80 636
rect 46 556 53 568
rect 73 556 80 568
rect 126 556 133 636
rect 188 627 195 654
rect 46 472 53 500
rect 73 472 80 500
rect 126 472 133 500
rect 188 472 195 611
rect 46 254 53 416
rect 73 254 80 416
rect 126 254 133 416
rect 46 196 53 224
rect 73 196 80 224
rect 126 196 133 224
rect 188 196 195 416
rect 216 409 223 654
rect 46 138 53 166
rect 73 138 80 166
rect 46 96 53 108
rect 73 96 80 108
rect 126 96 133 166
rect 188 139 195 166
rect 216 139 223 393
rect 188 101 195 109
rect 216 101 223 109
rect 46 57 53 66
rect 73 57 80 66
rect 126 57 133 66
<< ndiffusion >>
rect 43 224 46 254
rect 53 224 73 254
rect 80 224 126 254
rect 133 224 136 254
rect 43 166 46 196
rect 53 166 56 196
rect 70 166 73 196
rect 80 166 83 196
rect 97 166 126 196
rect 133 166 136 196
rect 185 166 188 196
rect 195 166 198 196
rect 43 108 46 138
rect 53 108 73 138
rect 80 108 83 138
rect 185 109 188 139
rect 195 109 198 139
rect 212 109 216 139
rect 223 109 226 139
rect 43 66 46 96
rect 53 66 56 96
rect 70 66 73 96
rect 80 66 83 96
rect 123 66 126 96
rect 133 66 136 96
<< pdiffusion >>
rect 43 636 46 692
rect 53 636 56 692
rect 70 636 73 692
rect 80 636 83 692
rect 123 636 126 692
rect 133 636 136 692
rect 185 654 188 710
rect 195 654 198 710
rect 212 654 216 710
rect 223 654 226 710
rect 43 568 46 624
rect 53 568 73 624
rect 80 568 83 624
rect 43 500 46 556
rect 53 500 56 556
rect 70 500 73 556
rect 80 500 83 556
rect 111 500 126 556
rect 133 500 136 556
rect 43 416 46 472
rect 53 416 73 472
rect 80 416 126 472
rect 133 416 136 472
rect 185 416 188 472
rect 195 416 198 472
<< ntransistor >>
rect 46 224 53 254
rect 73 224 80 254
rect 126 224 133 254
rect 46 166 53 196
rect 73 166 80 196
rect 126 166 133 196
rect 188 166 195 196
rect 46 108 53 138
rect 73 108 80 138
rect 188 109 195 139
rect 216 109 223 139
rect 46 66 53 96
rect 73 66 80 96
rect 126 66 133 96
<< ptransistor >>
rect 46 636 53 692
rect 73 636 80 692
rect 126 636 133 692
rect 188 654 195 710
rect 216 654 223 710
rect 46 568 53 624
rect 73 568 80 624
rect 46 500 53 556
rect 73 500 80 556
rect 126 500 133 556
rect 46 416 53 472
rect 73 416 80 472
rect 126 416 133 472
rect 188 416 195 472
<< polycontact >>
rect 37 701 53 717
rect 64 701 80 717
rect 117 701 133 717
rect 183 611 199 627
rect 212 393 228 409
rect 37 41 53 57
rect 64 41 80 57
rect 117 41 133 57
<< ndiffcontact >>
rect 29 224 43 254
rect 136 224 150 254
rect 29 166 43 196
rect 56 166 70 196
rect 83 166 97 196
rect 136 166 150 196
rect 171 166 185 196
rect 198 166 212 196
rect 29 108 43 138
rect 83 108 97 138
rect 171 109 185 139
rect 198 109 212 139
rect 226 109 240 139
rect 29 66 43 96
rect 56 66 70 96
rect 83 66 97 96
rect 109 66 123 96
rect 136 66 150 96
<< pdiffcontact >>
rect 29 636 43 692
rect 56 636 70 692
rect 83 636 97 692
rect 109 636 123 692
rect 136 636 150 692
rect 171 654 185 710
rect 198 654 212 710
rect 226 654 240 710
rect 29 568 43 624
rect 83 568 97 624
rect 29 500 43 556
rect 56 500 70 556
rect 83 500 111 556
rect 136 500 150 556
rect 29 416 43 472
rect 136 416 150 472
rect 171 416 185 472
rect 198 416 212 472
<< psubstratetap >>
rect 6 10 246 24
<< nsubstratetap >>
rect 6 734 246 748
<< metal1 >>
rect 0 748 252 752
rect 0 734 6 748
rect 246 734 252 748
rect 0 728 252 734
rect 9 692 26 728
rect 90 692 100 728
rect 198 710 212 728
rect 9 636 29 692
rect 97 636 100 692
rect 9 556 20 636
rect 136 624 150 636
rect 97 614 112 624
rect 130 614 183 624
rect 9 541 29 556
rect 9 536 23 541
rect 56 491 70 500
rect 136 491 150 500
rect 56 481 150 491
rect 136 472 150 481
rect 150 416 171 472
rect 29 407 43 416
rect 198 407 212 416
rect 29 397 154 407
rect 172 397 212 407
rect 0 370 252 380
rect 0 351 252 361
rect 0 307 252 317
rect 0 288 252 298
rect 0 263 252 273
rect 29 196 43 224
rect 56 205 208 215
rect 56 196 70 205
rect 136 196 150 205
rect 198 196 208 205
rect 29 157 43 166
rect 83 157 97 166
rect 29 147 97 157
rect 29 138 43 147
rect 29 96 43 108
rect 16 66 29 96
rect 97 66 100 96
rect 16 30 26 66
rect 90 30 100 66
rect 198 30 212 109
rect 0 24 252 30
rect 0 10 6 24
rect 246 10 252 24
rect 0 6 252 10
<< m2contact >>
rect 35 717 53 719
rect 35 701 37 717
rect 37 701 53 717
rect 63 717 81 719
rect 63 701 64 717
rect 64 701 80 717
rect 80 701 81 717
rect 115 717 133 719
rect 115 701 117 717
rect 117 701 133 717
rect 54 636 56 654
rect 56 636 70 654
rect 70 636 72 654
rect 109 636 123 654
rect 123 636 127 654
rect 165 670 171 688
rect 171 670 183 688
rect 228 670 240 688
rect 240 670 246 688
rect 29 606 43 624
rect 43 606 47 624
rect 112 606 130 624
rect 23 521 29 541
rect 29 521 43 541
rect 87 519 107 539
rect 154 389 172 407
rect 136 229 150 247
rect 150 229 154 247
rect 167 171 171 189
rect 171 171 185 189
rect 82 118 83 136
rect 83 118 97 136
rect 97 118 100 136
rect 167 119 171 137
rect 171 119 185 137
rect 226 119 240 137
rect 240 119 244 137
rect 54 78 56 96
rect 56 78 70 96
rect 70 78 72 96
rect 109 78 123 96
rect 123 78 127 96
rect 137 78 150 96
rect 150 78 155 96
rect 35 41 37 57
rect 37 41 53 57
rect 35 39 53 41
rect 63 41 64 57
rect 64 41 80 57
rect 80 41 81 57
rect 63 39 81 41
rect 115 41 117 57
rect 117 41 133 57
rect 115 39 133 41
<< metal2 >>
rect 28 719 40 758
rect 56 745 68 758
rect 56 733 75 745
rect 63 719 75 733
rect 112 719 124 758
rect 196 726 208 758
rect 28 701 35 719
rect 112 701 115 719
rect 182 713 208 726
rect 224 725 236 758
rect 224 713 244 725
rect 182 688 194 713
rect 232 688 244 713
rect 183 670 194 688
rect 72 636 109 648
rect 35 624 66 636
rect 43 523 87 535
rect 117 486 129 606
rect 110 474 129 486
rect 110 136 122 474
rect 160 247 172 389
rect 154 229 172 247
rect 160 189 172 229
rect 182 228 194 670
rect 182 216 211 228
rect 160 171 167 189
rect 199 160 211 216
rect 182 148 211 160
rect 182 137 194 148
rect 232 137 244 670
rect 100 130 122 136
rect 100 118 149 130
rect 185 119 194 137
rect 60 96 121 108
rect 137 96 149 118
rect 28 39 35 57
rect 28 0 40 39
rect 63 27 81 39
rect 56 15 81 27
rect 112 39 115 57
rect 56 0 68 15
rect 112 0 124 39
rect 182 38 194 119
rect 182 26 208 38
rect 232 37 244 119
rect 196 0 208 26
rect 224 25 244 37
rect 224 0 236 25
<< labels >>
rlabel metal1 252 6 252 30 7 GND!
rlabel metal1 0 6 0 30 3 GND!
rlabel metal2 28 0 40 0 1 A
rlabel metal2 56 0 68 0 1 B
rlabel metal2 112 0 124 0 1 Cin
rlabel metal2 196 0 208 0 1 Cout
rlabel metal2 224 0 236 0 1 S
rlabel metal1 0 263 0 273 3 nReset
rlabel metal1 0 288 0 298 3 Clock
rlabel metal1 0 307 0 317 3 Test
rlabel metal1 0 351 0 361 3 Scan
rlabel metal1 0 370 0 380 3 ScanReturn
rlabel metal1 252 370 252 380 7 ScanReturn
rlabel metal1 252 351 252 361 7 Scan
rlabel metal1 252 307 252 317 7 Test
rlabel metal1 252 288 252 298 7 Clock
rlabel metal1 252 263 252 273 7 nReset
rlabel metal1 0 728 0 752 3 Vdd!
rlabel metal1 252 728 252 752 7 Vdd!
rlabel metal2 28 758 40 758 5 A
rlabel metal2 196 758 208 758 5 Cout
rlabel metal2 224 758 236 758 5 S
rlabel metal2 112 758 124 758 5 Cin
rlabel metal2 56 758 68 758 5 B
<< end >>
