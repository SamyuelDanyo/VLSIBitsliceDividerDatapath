magic
tech c35b4
timestamp 1544089383
<< pimplant >>
rect 1165 334 1316 727
<< nimplant >>
rect 1165 31 1316 281
<< nwell >>
rect 327 446 1316 752
rect 437 351 1316 446
rect 688 334 1316 351
<< polysilicon >>
rect 373 719 380 727
rect 402 719 409 727
rect 455 719 462 727
rect 482 719 489 727
rect 535 719 542 727
rect 562 719 569 727
rect 615 719 622 727
rect 668 719 675 727
rect 695 719 702 727
rect 749 719 756 727
rect 776 719 783 727
rect 830 719 837 727
rect 857 719 864 727
rect 911 719 918 727
rect 938 719 945 727
rect 965 719 972 727
rect 992 719 999 727
rect 1045 719 1052 727
rect 1072 719 1079 727
rect 1099 719 1106 727
rect 1126 719 1133 727
rect 1179 719 1186 727
rect 1206 719 1213 727
rect 1233 719 1240 727
rect 1260 719 1267 727
rect 373 330 380 663
rect 373 314 377 330
rect 373 69 380 314
rect 402 276 409 653
rect 402 59 409 260
rect 455 248 462 653
rect 455 59 462 232
rect 482 214 489 653
rect 535 439 542 540
rect 562 465 569 540
rect 615 496 622 540
rect 482 59 489 198
rect 535 93 542 423
rect 562 93 569 449
rect 615 93 622 480
rect 668 408 675 478
rect 695 403 702 478
rect 684 396 702 403
rect 668 112 675 392
rect 695 112 702 396
rect 749 435 756 478
rect 776 430 783 478
rect 765 423 783 430
rect 749 112 756 419
rect 776 112 783 423
rect 830 460 837 478
rect 857 455 864 478
rect 846 448 864 455
rect 830 112 837 444
rect 857 112 864 448
rect 911 380 918 389
rect 938 375 945 389
rect 965 375 972 389
rect 992 375 999 389
rect 927 368 999 375
rect 911 139 918 364
rect 938 139 945 368
rect 965 139 972 368
rect 992 139 999 368
rect 1045 360 1052 389
rect 1072 353 1079 389
rect 1099 353 1106 389
rect 1126 353 1133 389
rect 1052 346 1133 353
rect 1045 139 1052 344
rect 1072 139 1079 346
rect 1099 139 1106 346
rect 1126 139 1133 346
rect 1179 341 1186 389
rect 1177 334 1186 341
rect 1206 334 1213 389
rect 1233 334 1240 389
rect 1260 334 1267 389
rect 1177 327 1267 334
rect 1177 325 1186 327
rect 1179 139 1186 325
rect 1206 139 1213 327
rect 1233 139 1240 327
rect 1260 139 1267 327
rect 373 31 380 39
rect 402 31 409 39
rect 455 31 462 39
rect 482 31 489 39
rect 535 31 542 39
rect 562 31 569 39
rect 615 31 622 39
rect 668 31 675 39
rect 695 31 702 39
rect 749 31 756 39
rect 776 31 783 39
rect 830 31 837 39
rect 857 31 864 39
rect 911 31 918 39
rect 938 31 945 39
rect 965 31 972 39
rect 992 31 999 39
rect 1045 31 1052 39
rect 1072 31 1079 39
rect 1099 31 1106 39
rect 1126 31 1133 39
rect 1179 31 1186 39
rect 1206 31 1213 39
rect 1233 31 1240 39
rect 1260 31 1267 39
<< ndiffusion >>
rect 370 39 373 69
rect 380 39 384 69
rect 398 39 402 59
rect 409 39 412 59
rect 452 39 455 59
rect 462 39 465 59
rect 479 39 482 59
rect 489 39 492 59
rect 532 39 535 93
rect 542 39 545 93
rect 559 39 562 93
rect 569 39 572 93
rect 612 39 615 93
rect 622 39 625 93
rect 665 39 668 112
rect 675 39 678 112
rect 692 39 695 112
rect 702 39 705 112
rect 746 39 749 112
rect 756 39 759 112
rect 773 39 776 112
rect 783 39 786 112
rect 827 39 830 112
rect 837 39 840 112
rect 854 39 857 112
rect 864 39 867 112
rect 908 39 911 139
rect 918 39 921 139
rect 935 39 938 139
rect 945 39 948 139
rect 962 39 965 139
rect 972 39 975 139
rect 989 39 992 139
rect 999 39 1002 139
rect 1042 39 1045 139
rect 1052 39 1055 139
rect 1069 39 1072 139
rect 1079 39 1082 139
rect 1096 39 1099 139
rect 1106 39 1109 139
rect 1123 39 1126 139
rect 1133 39 1136 139
rect 1176 39 1179 139
rect 1186 39 1189 139
rect 1203 39 1206 139
rect 1213 39 1216 139
rect 1230 39 1233 139
rect 1240 39 1243 139
rect 1257 39 1260 139
rect 1267 39 1270 139
<< pdiffusion >>
rect 370 663 373 719
rect 380 663 384 719
rect 398 653 402 719
rect 409 653 412 719
rect 452 653 455 719
rect 462 653 465 719
rect 479 653 482 719
rect 489 653 492 719
rect 532 540 535 719
rect 542 540 545 719
rect 559 540 562 719
rect 569 540 572 719
rect 612 540 615 719
rect 622 540 625 719
rect 665 478 668 719
rect 675 478 678 719
rect 692 478 695 719
rect 702 478 705 719
rect 746 478 749 719
rect 756 478 759 719
rect 773 478 776 719
rect 783 478 786 719
rect 827 478 830 719
rect 837 478 840 719
rect 854 478 857 719
rect 864 478 867 719
rect 908 389 911 719
rect 918 389 921 719
rect 935 389 938 719
rect 945 389 948 719
rect 962 389 965 719
rect 972 389 975 719
rect 989 389 992 719
rect 999 389 1002 719
rect 1042 389 1045 719
rect 1052 389 1055 719
rect 1069 389 1072 719
rect 1079 389 1082 719
rect 1096 389 1099 719
rect 1106 389 1109 719
rect 1123 389 1126 719
rect 1133 389 1136 719
rect 1176 389 1179 719
rect 1186 389 1189 719
rect 1203 389 1206 719
rect 1213 389 1216 719
rect 1230 389 1233 719
rect 1240 389 1243 719
rect 1257 389 1260 719
rect 1267 389 1270 719
<< ntransistor >>
rect 373 39 380 69
rect 402 39 409 59
rect 455 39 462 59
rect 482 39 489 59
rect 535 39 542 93
rect 562 39 569 93
rect 615 39 622 93
rect 668 39 675 112
rect 695 39 702 112
rect 749 39 756 112
rect 776 39 783 112
rect 830 39 837 112
rect 857 39 864 112
rect 911 39 918 139
rect 938 39 945 139
rect 965 39 972 139
rect 992 39 999 139
rect 1045 39 1052 139
rect 1072 39 1079 139
rect 1099 39 1106 139
rect 1126 39 1133 139
rect 1179 39 1186 139
rect 1206 39 1213 139
rect 1233 39 1240 139
rect 1260 39 1267 139
<< ptransistor >>
rect 373 663 380 719
rect 402 653 409 719
rect 455 653 462 719
rect 482 653 489 719
rect 535 540 542 719
rect 562 540 569 719
rect 615 540 622 719
rect 668 478 675 719
rect 695 478 702 719
rect 749 478 756 719
rect 776 478 783 719
rect 830 478 837 719
rect 857 478 864 719
rect 911 389 918 719
rect 938 389 945 719
rect 965 389 972 719
rect 992 389 999 719
rect 1045 389 1052 719
rect 1072 389 1079 719
rect 1099 389 1106 719
rect 1126 389 1133 719
rect 1179 389 1186 719
rect 1206 389 1213 719
rect 1233 389 1240 719
rect 1260 389 1267 719
<< polycontact >>
rect 0 12 239 680
rect 377 314 393 330
rect 393 260 409 276
rect 446 232 462 248
rect 606 480 622 496
rect 553 449 569 465
rect 526 423 542 439
rect 473 198 489 214
rect 668 392 684 408
rect 749 419 765 435
rect 830 444 846 460
rect 911 364 927 380
rect 1036 344 1052 360
rect 1161 325 1177 341
<< ndiffcontact >>
rect 356 39 370 69
rect 384 39 398 69
rect 412 39 426 59
rect 438 39 452 59
rect 465 39 479 59
rect 492 39 506 59
rect 518 39 532 93
rect 545 39 559 93
rect 572 39 586 93
rect 598 39 612 93
rect 625 39 639 93
rect 651 39 665 112
rect 678 39 692 112
rect 705 39 719 112
rect 732 39 746 112
rect 759 39 773 112
rect 786 39 800 112
rect 813 39 827 112
rect 840 39 854 112
rect 867 39 881 112
rect 894 39 908 139
rect 921 39 935 139
rect 948 39 962 139
rect 975 39 989 139
rect 1002 39 1016 139
rect 1028 39 1042 139
rect 1055 39 1069 139
rect 1082 39 1096 139
rect 1109 39 1123 139
rect 1136 39 1150 139
rect 1162 39 1176 139
rect 1189 39 1203 139
rect 1216 39 1230 139
rect 1243 39 1257 139
rect 1270 39 1284 139
<< pdiffcontact >>
rect 356 663 370 719
rect 384 653 398 719
rect 412 653 426 719
rect 438 653 452 719
rect 465 653 479 719
rect 492 653 506 719
rect 518 540 532 719
rect 545 540 559 719
rect 572 540 586 719
rect 598 540 612 719
rect 625 540 639 719
rect 651 478 665 719
rect 678 478 692 719
rect 705 478 719 719
rect 732 478 746 719
rect 759 478 773 719
rect 786 478 800 719
rect 813 478 827 719
rect 840 478 854 719
rect 867 478 881 719
rect 894 389 908 719
rect 921 389 935 719
rect 948 389 962 719
rect 975 389 989 719
rect 1002 389 1016 719
rect 1028 389 1042 719
rect 1055 389 1069 719
rect 1082 389 1096 719
rect 1109 389 1123 719
rect 1136 389 1150 719
rect 1162 389 1176 719
rect 1189 389 1203 719
rect 1216 389 1230 719
rect 1243 389 1257 719
rect 1270 389 1284 719
<< psubstratetap >>
rect 337 10 1310 24
<< nsubstratetap >>
rect 332 734 1310 748
<< metal1 >>
rect 240 748 1316 752
rect 240 734 332 748
rect 1310 734 1316 748
rect 240 728 1316 734
rect 384 719 398 728
rect 465 719 479 728
rect 545 719 559 728
rect 598 719 612 728
rect 678 719 692 728
rect 759 719 773 728
rect 840 719 854 728
rect 921 719 935 728
rect 975 719 989 728
rect 1055 719 1069 728
rect 1109 719 1123 728
rect 1189 719 1203 728
rect 1243 719 1257 728
rect 357 374 369 663
rect 414 611 424 653
rect 440 640 450 653
rect 494 640 504 653
rect 520 531 530 540
rect 574 531 584 540
rect 627 530 637 540
rect 504 483 606 493
rect 457 451 553 461
rect 643 447 830 457
rect 426 426 526 436
rect 591 422 749 432
rect 536 395 668 405
rect 722 370 911 380
rect 1187 370 1316 380
rect 804 345 1036 355
rect 274 317 350 327
rect 393 315 843 325
rect 879 325 1161 335
rect 1187 316 1197 370
rect 833 309 843 315
rect 888 309 1197 316
rect 833 306 1197 309
rect 1207 351 1316 361
rect 274 295 824 305
rect 833 299 898 306
rect 1207 297 1217 351
rect 814 290 824 295
rect 907 290 1217 297
rect 814 287 1217 290
rect 1226 307 1316 317
rect 814 280 917 287
rect 1226 278 1236 307
rect 296 266 393 276
rect 1016 268 1236 278
rect 1245 288 1316 298
rect 325 237 446 247
rect 347 201 473 211
rect 359 69 369 128
rect 414 59 424 110
rect 520 93 530 119
rect 574 93 584 119
rect 653 112 663 141
rect 707 112 717 176
rect 734 112 744 148
rect 788 112 798 131
rect 815 112 825 163
rect 869 112 879 154
rect 896 139 906 185
rect 951 139 961 185
rect 1004 139 1014 260
rect 1245 259 1255 288
rect 1150 249 1255 259
rect 1285 263 1316 273
rect 1030 139 1040 199
rect 1083 139 1093 159
rect 1138 139 1148 241
rect 1164 139 1174 198
rect 1218 139 1228 198
rect 1273 139 1283 255
rect 627 93 637 108
rect 441 59 451 77
rect 494 59 504 68
rect 384 30 398 39
rect 465 30 479 39
rect 545 30 559 39
rect 598 30 612 39
rect 678 30 692 39
rect 759 30 773 39
rect 840 30 854 39
rect 921 30 935 39
rect 975 30 989 39
rect 1055 30 1069 39
rect 1109 30 1123 39
rect 1189 30 1203 39
rect 1243 30 1257 39
rect 276 24 1316 30
rect 276 10 337 24
rect 1310 10 1316 24
rect 276 6 1316 10
<< m2contact >>
rect 0 728 240 752
rect 0 12 239 680
rect 436 622 454 640
rect 491 622 509 640
rect 411 593 429 611
rect 514 513 532 531
rect 571 513 589 531
rect 619 512 637 530
rect 647 508 651 526
rect 651 508 665 526
rect 486 478 504 496
rect 728 508 732 526
rect 732 508 746 526
rect 705 478 719 496
rect 719 478 723 496
rect 809 508 813 526
rect 813 508 827 526
rect 786 478 800 496
rect 800 478 804 496
rect 866 478 867 496
rect 867 478 881 496
rect 881 478 884 496
rect 439 447 457 465
rect 625 443 643 461
rect 408 422 426 440
rect 573 418 591 436
rect 518 391 536 409
rect 890 389 894 407
rect 894 389 908 407
rect 1025 417 1028 435
rect 1028 417 1042 435
rect 1042 417 1043 435
rect 1159 417 1162 435
rect 1162 417 1176 435
rect 1176 417 1177 435
rect 1135 389 1136 407
rect 1136 389 1150 407
rect 1150 389 1153 407
rect 1215 389 1216 407
rect 1216 389 1230 407
rect 1230 389 1233 407
rect 1269 389 1270 407
rect 1270 389 1284 407
rect 1284 389 1287 407
rect 356 356 374 374
rect 704 366 722 384
rect 946 371 964 389
rect 1001 371 1019 389
rect 1080 371 1098 389
rect 786 343 804 361
rect 256 315 274 333
rect 350 314 368 332
rect 861 318 879 336
rect 256 287 274 305
rect 278 258 296 276
rect 998 260 1016 278
rect 307 229 325 247
rect 329 195 347 213
rect 705 176 723 194
rect 892 185 910 203
rect 946 185 964 203
rect 357 128 375 146
rect 648 141 666 159
rect 411 110 429 128
rect 516 119 534 137
rect 571 119 589 137
rect 436 77 454 95
rect 624 108 642 126
rect 729 148 747 166
rect 810 163 828 181
rect 786 131 804 149
rect 867 154 885 172
rect 1132 241 1150 259
rect 1267 255 1285 273
rect 1027 199 1045 217
rect 1079 159 1097 177
rect 1161 198 1179 216
rect 1214 198 1232 216
rect 490 68 508 86
<< metal2 >>
rect 0 752 240 758
rect 0 680 240 728
rect 239 12 240 680
rect 280 651 292 758
rect 262 639 292 651
rect 262 333 274 639
rect 308 629 320 758
rect 284 617 320 629
rect 256 52 268 287
rect 284 276 296 617
rect 336 607 348 758
rect 306 595 348 607
rect 306 276 318 595
rect 364 585 376 758
rect 330 573 376 585
rect 330 354 342 573
rect 414 440 426 593
rect 328 342 342 354
rect 328 298 340 342
rect 357 332 369 356
rect 368 314 369 332
rect 328 286 347 298
rect 306 264 319 276
rect 284 74 296 258
rect 307 247 319 264
rect 307 96 319 229
rect 335 213 347 286
rect 335 118 347 195
rect 357 146 369 314
rect 414 128 426 422
rect 439 465 451 622
rect 492 496 504 622
rect 335 106 376 118
rect 307 84 348 96
rect 284 62 320 74
rect 256 40 292 52
rect 0 0 240 12
rect 280 0 292 40
rect 308 0 320 62
rect 336 0 348 84
rect 364 0 376 106
rect 439 95 451 447
rect 492 86 504 478
rect 518 409 530 513
rect 573 436 585 513
rect 625 461 637 512
rect 653 444 665 508
rect 705 444 717 478
rect 518 137 530 391
rect 573 137 585 418
rect 625 126 637 443
rect 653 432 717 444
rect 653 159 665 432
rect 705 384 717 432
rect 734 447 746 508
rect 786 447 798 478
rect 734 435 798 447
rect 705 194 717 366
rect 734 166 746 435
rect 786 361 798 435
rect 815 444 827 508
rect 867 444 879 478
rect 815 432 879 444
rect 786 149 798 343
rect 815 181 827 432
rect 867 336 879 432
rect 867 172 879 318
rect 895 377 907 389
rect 895 371 946 377
rect 964 371 1001 377
rect 1029 377 1041 417
rect 1029 371 1080 377
rect 1138 377 1150 389
rect 1098 371 1150 377
rect 895 365 1016 371
rect 895 203 907 365
rect 949 203 961 365
rect 1004 278 1016 365
rect 1029 365 1150 371
rect 1029 217 1041 365
rect 1083 177 1095 365
rect 1138 259 1150 365
rect 1163 378 1175 417
rect 1219 378 1231 389
rect 1272 378 1284 389
rect 1163 366 1284 378
rect 1163 216 1175 366
rect 1219 216 1231 366
rect 1272 273 1284 366
<< labels >>
rlabel metal1 1316 370 1316 380 7 nSDO
rlabel metal1 1316 6 1316 30 7 GND!
rlabel metal1 1316 728 1316 752 7 Vdd!
rlabel metal1 1316 351 1316 361 7 SDI
rlabel metal1 1316 263 1316 273 7 nResetOut
rlabel metal1 1316 288 1316 298 7 ClockOut
rlabel metal1 1316 307 1316 317 7 TestOut
rlabel metal2 364 758 376 758 5 nReset
rlabel metal2 336 758 348 758 5 Clock
rlabel metal2 308 758 320 758 5 Test
rlabel metal2 280 758 292 758 5 SDO
rlabel metal2 0 758 240 758 5 Vdd!
rlabel metal2 0 0 240 0 1 Vdd!
rlabel metal2 364 0 376 0 1 nReset
rlabel metal2 336 0 348 0 1 Clock
rlabel metal2 308 0 320 0 1 Test
rlabel metal2 280 0 292 0 1 SDI
<< end >>
