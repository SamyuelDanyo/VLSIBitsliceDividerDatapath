magic
tech c35b4
timestamp 1543772215
<< pimplant >>
rect 0 334 588 727
<< nimplant >>
rect 0 31 588 281
<< nwell >>
rect 0 334 588 752
<< polysilicon >>
rect 23 715 30 724
rect 51 715 58 724
rect 23 631 30 659
rect 51 631 58 659
rect 78 631 85 724
rect 105 631 112 724
rect 191 624 198 727
rect 219 692 226 727
rect 247 692 254 727
rect 300 717 307 727
rect 300 701 306 717
rect 300 692 307 701
rect 333 692 340 727
rect 372 692 379 727
rect 425 692 432 727
rect 219 624 226 636
rect 23 323 30 575
rect 23 131 30 307
rect 51 131 58 575
rect 78 526 85 575
rect 78 131 85 508
rect 105 361 112 575
rect 247 571 254 636
rect 300 624 307 636
rect 191 540 198 568
rect 219 555 226 568
rect 247 564 279 571
rect 219 548 251 555
rect 244 540 251 548
rect 105 131 112 345
rect 191 298 198 484
rect 244 374 251 484
rect 219 367 251 374
rect 191 235 198 282
rect 219 279 226 367
rect 272 358 279 564
rect 300 555 307 568
rect 333 555 340 636
rect 372 624 379 636
rect 425 624 432 636
rect 372 560 379 568
rect 247 351 279 358
rect 288 548 307 555
rect 316 548 340 555
rect 369 553 379 560
rect 425 555 432 568
rect 458 567 465 727
rect 247 342 254 351
rect 247 303 254 326
rect 247 296 279 303
rect 219 247 226 263
rect 219 240 251 247
rect 244 235 251 240
rect 191 155 198 205
rect 244 200 251 205
rect 219 193 251 200
rect 219 155 226 193
rect 23 73 30 101
rect 51 73 58 101
rect 23 34 30 43
rect 51 34 58 43
rect 78 34 85 101
rect 105 34 112 101
rect 191 31 198 125
rect 219 113 226 125
rect 272 113 279 296
rect 288 166 295 548
rect 316 540 323 548
rect 369 540 376 553
rect 422 548 432 555
rect 449 549 458 556
rect 422 540 429 548
rect 449 540 456 549
rect 502 540 509 727
rect 316 358 323 484
rect 369 358 376 484
rect 422 475 429 484
rect 422 468 424 475
rect 429 358 436 457
rect 316 351 328 358
rect 369 351 386 358
rect 429 351 439 358
rect 321 235 328 351
rect 379 235 386 351
rect 432 235 439 351
rect 449 260 456 484
rect 502 475 509 484
rect 448 235 455 244
rect 501 235 508 459
rect 321 182 328 205
rect 321 175 366 182
rect 288 159 332 166
rect 325 155 332 159
rect 325 113 332 125
rect 359 85 366 175
rect 379 171 386 205
rect 432 180 439 205
rect 448 201 455 205
rect 448 194 490 201
rect 379 164 409 171
rect 448 164 462 171
rect 402 155 409 164
rect 455 155 462 164
rect 402 113 409 125
rect 455 113 462 125
rect 219 31 226 83
rect 272 31 279 83
rect 325 74 332 83
rect 325 31 332 58
rect 361 31 368 67
rect 402 31 409 83
rect 455 31 462 83
rect 483 74 490 194
rect 501 102 508 205
rect 483 31 490 56
rect 501 31 508 84
<< ndiffusion >>
rect 188 205 191 235
rect 198 205 201 235
rect 241 205 244 235
rect 251 205 254 235
rect 20 101 23 131
rect 30 101 33 131
rect 47 101 51 131
rect 58 101 78 131
rect 85 101 88 131
rect 102 101 105 131
rect 112 101 115 131
rect 188 125 191 155
rect 198 125 219 155
rect 226 125 229 155
rect 20 43 23 73
rect 30 43 33 73
rect 318 205 321 235
rect 328 205 336 235
rect 376 205 379 235
rect 386 205 389 235
rect 429 205 432 235
rect 439 205 448 235
rect 455 205 458 235
rect 498 205 501 235
rect 508 205 511 235
rect 322 125 325 155
rect 332 125 335 155
rect 216 83 219 113
rect 226 83 229 113
rect 269 83 272 113
rect 279 83 282 113
rect 322 83 325 113
rect 332 83 335 113
rect 452 125 455 155
rect 462 125 465 155
rect 399 83 402 113
rect 409 83 412 113
rect 452 83 455 113
rect 462 83 465 113
<< pdiffusion >>
rect 20 659 23 715
rect 30 659 33 715
rect 20 575 23 631
rect 30 575 33 631
rect 47 575 51 631
rect 58 575 61 631
rect 75 575 78 631
rect 85 575 88 631
rect 102 575 105 631
rect 112 575 115 631
rect 216 636 219 692
rect 226 636 229 692
rect 243 636 247 692
rect 254 636 257 692
rect 297 636 300 692
rect 307 636 310 692
rect 369 636 372 692
rect 379 636 382 692
rect 422 636 425 692
rect 432 636 435 692
rect 188 568 191 624
rect 198 568 201 624
rect 216 568 219 624
rect 226 568 229 624
rect 297 568 300 624
rect 307 568 310 624
rect 188 484 191 540
rect 198 484 201 540
rect 241 484 244 540
rect 251 484 254 540
rect 422 568 425 624
rect 432 568 435 624
rect 313 484 316 540
rect 323 484 326 540
rect 366 484 369 540
rect 376 484 379 540
rect 419 484 422 540
rect 429 484 432 540
rect 446 484 449 540
rect 456 484 459 540
rect 499 484 502 540
rect 509 484 512 540
<< ntransistor >>
rect 191 205 198 235
rect 244 205 251 235
rect 23 101 30 131
rect 51 101 58 131
rect 78 101 85 131
rect 105 101 112 131
rect 191 125 198 155
rect 219 125 226 155
rect 23 43 30 73
rect 321 205 328 235
rect 379 205 386 235
rect 432 205 439 235
rect 448 205 455 235
rect 501 205 508 235
rect 325 125 332 155
rect 219 83 226 113
rect 272 83 279 113
rect 325 83 332 113
rect 455 125 462 155
rect 402 83 409 113
rect 455 83 462 113
<< ptransistor >>
rect 23 659 30 715
rect 23 575 30 631
rect 51 575 58 631
rect 78 575 85 631
rect 105 575 112 631
rect 219 636 226 692
rect 247 636 254 692
rect 300 636 307 692
rect 372 636 379 692
rect 425 636 432 692
rect 191 568 198 624
rect 219 568 226 624
rect 300 568 307 624
rect 191 484 198 540
rect 244 484 251 540
rect 425 568 432 624
rect 316 484 323 540
rect 369 484 376 540
rect 422 484 429 540
rect 449 484 456 540
rect 502 484 509 540
<< polycontact >>
rect 51 659 67 715
rect 306 701 322 717
rect 328 636 344 692
rect 22 307 38 323
rect 78 508 96 526
rect 105 345 121 361
rect 187 282 203 298
rect 372 568 388 624
rect 242 326 258 342
rect 215 263 231 279
rect 51 43 67 73
rect 458 549 474 567
rect 424 457 440 475
rect 499 459 515 475
rect 448 244 464 260
rect 432 164 448 180
rect 393 125 409 155
rect 322 58 338 74
rect 359 67 375 85
rect 499 84 515 102
rect 474 56 490 74
<< ndiffcontact >>
rect 174 205 188 235
rect 201 205 215 235
rect 227 205 241 235
rect 254 205 268 235
rect 6 101 20 131
rect 33 101 47 131
rect 88 101 102 131
rect 115 101 129 131
rect 174 125 188 155
rect 229 125 243 155
rect 6 43 20 73
rect 33 43 47 73
rect 304 205 318 235
rect 336 205 350 235
rect 362 205 376 235
rect 389 205 403 235
rect 415 205 429 235
rect 458 205 472 235
rect 484 205 498 235
rect 511 205 525 235
rect 308 125 322 155
rect 335 125 349 155
rect 202 83 216 113
rect 229 83 243 113
rect 255 83 269 113
rect 282 83 296 113
rect 308 83 322 113
rect 335 83 349 113
rect 438 125 452 155
rect 465 125 479 155
rect 385 83 399 113
rect 412 83 426 113
rect 438 83 452 113
rect 465 83 479 113
<< pdiffcontact >>
rect 6 659 20 715
rect 33 659 47 715
rect 6 575 20 631
rect 33 575 47 631
rect 61 575 75 631
rect 88 575 102 631
rect 115 575 129 631
rect 202 636 216 692
rect 229 636 243 692
rect 257 636 271 692
rect 283 636 297 692
rect 310 636 324 692
rect 355 636 369 692
rect 382 636 396 692
rect 408 636 422 692
rect 435 636 449 692
rect 174 568 188 624
rect 201 568 216 624
rect 229 568 243 624
rect 283 568 297 624
rect 310 568 324 624
rect 174 484 188 540
rect 201 484 215 540
rect 227 484 241 540
rect 254 484 268 540
rect 408 568 422 624
rect 435 568 449 624
rect 299 484 313 540
rect 326 484 340 540
rect 352 484 366 540
rect 379 484 393 540
rect 405 484 419 540
rect 432 484 446 540
rect 459 484 473 540
rect 485 484 499 540
rect 512 484 526 540
<< psubstratetap >>
rect 6 10 582 24
<< nsubstratetap >>
rect 6 734 582 748
<< metal1 >>
rect 0 748 588 752
rect 0 734 6 748
rect 582 734 588 748
rect 0 728 588 734
rect 6 715 20 728
rect 47 659 51 715
rect 6 631 20 659
rect 35 640 100 650
rect 35 631 45 640
rect 90 631 100 640
rect 115 631 129 728
rect 174 624 188 728
rect 229 692 243 728
rect 283 692 297 728
rect 324 701 369 717
rect 355 692 369 701
rect 324 636 328 692
rect 382 692 396 728
rect 435 692 449 728
rect 63 566 73 575
rect 324 620 372 624
rect 326 602 372 620
rect 324 568 372 602
rect 388 568 408 624
rect 63 556 124 566
rect 174 540 188 568
rect 379 549 458 559
rect 474 549 499 559
rect 379 540 393 549
rect 485 540 499 549
rect 254 475 268 484
rect 405 475 415 484
rect 459 475 473 484
rect 254 465 415 475
rect 459 459 499 475
rect 0 370 588 380
rect 0 351 105 361
rect 168 351 532 361
rect 550 351 588 361
rect 148 329 242 339
rect 0 307 22 317
rect 38 307 588 317
rect 0 288 187 298
rect 203 288 588 298
rect 0 263 215 273
rect 400 273 498 279
rect 231 269 588 273
rect 231 263 410 269
rect 488 263 588 269
rect 201 244 318 254
rect 464 244 498 254
rect 201 235 215 244
rect 304 235 318 244
rect 484 235 498 244
rect 35 159 124 170
rect 35 131 45 159
rect 174 155 188 205
rect 336 174 350 205
rect 458 196 472 205
rect 458 186 515 196
rect 336 164 432 174
rect 63 140 127 150
rect 8 92 18 101
rect 63 92 73 140
rect 116 131 127 140
rect 8 82 73 92
rect 243 125 308 155
rect 409 125 438 155
rect 174 113 188 125
rect 47 43 51 73
rect 6 30 20 43
rect 88 30 102 101
rect 174 83 202 113
rect 174 30 188 83
rect 255 49 269 83
rect 282 74 296 83
rect 282 58 322 74
rect 385 49 399 83
rect 255 39 399 49
rect 499 102 515 186
rect 412 30 426 83
rect 515 84 560 102
rect 490 56 532 74
rect 0 24 588 30
rect 0 10 6 24
rect 582 10 588 24
rect 0 6 588 10
<< m2contact >>
rect 306 717 324 719
rect 306 701 322 717
rect 322 701 324 717
rect 200 636 202 654
rect 202 636 216 654
rect 216 636 218 654
rect 255 674 257 692
rect 257 674 271 692
rect 271 674 273 692
rect 306 636 310 654
rect 310 636 324 654
rect 406 636 408 654
rect 408 636 422 654
rect 422 636 424 654
rect 200 602 201 620
rect 201 602 216 620
rect 216 602 218 620
rect 174 574 188 592
rect 188 574 192 592
rect 308 602 310 620
rect 310 602 324 620
rect 324 602 326 620
rect 227 574 229 592
rect 229 574 243 592
rect 243 574 245 592
rect 281 574 283 592
rect 283 574 297 592
rect 297 574 299 592
rect 431 574 435 592
rect 435 574 449 592
rect 124 548 142 566
rect 78 508 96 526
rect 174 522 188 540
rect 188 522 192 540
rect 225 522 227 540
rect 227 522 241 540
rect 241 522 243 540
rect 199 494 201 512
rect 201 494 215 512
rect 215 494 217 512
rect 297 522 299 540
rect 299 522 313 540
rect 313 522 315 540
rect 350 522 352 540
rect 352 522 366 540
rect 366 522 368 540
rect 324 494 326 512
rect 326 494 340 512
rect 340 494 342 512
rect 430 522 432 540
rect 432 522 446 540
rect 446 522 448 540
rect 403 494 405 512
rect 405 494 419 512
rect 419 494 421 512
rect 458 494 459 512
rect 459 494 473 512
rect 473 494 476 512
rect 510 522 512 540
rect 512 522 526 540
rect 526 522 528 540
rect 424 457 440 475
rect 440 457 442 475
rect 130 329 148 347
rect 532 343 550 361
rect 174 217 188 235
rect 188 217 192 235
rect 225 217 227 235
rect 227 217 241 235
rect 241 217 243 235
rect 252 205 254 207
rect 254 205 268 207
rect 268 205 270 207
rect 359 217 362 235
rect 362 217 376 235
rect 376 217 377 235
rect 387 217 389 235
rect 389 217 403 235
rect 403 217 405 235
rect 413 205 415 207
rect 415 205 429 207
rect 429 205 431 207
rect 124 159 142 177
rect 252 189 270 205
rect 413 189 431 205
rect 509 217 511 235
rect 511 217 525 235
rect 525 217 527 235
rect 333 137 335 155
rect 335 137 349 155
rect 349 137 351 155
rect 463 137 465 155
rect 465 137 479 155
rect 479 137 481 155
rect 226 95 229 113
rect 229 95 243 113
rect 243 95 244 113
rect 305 95 308 113
rect 308 95 322 113
rect 322 95 323 113
rect 333 95 335 113
rect 335 95 349 113
rect 349 95 351 113
rect 358 67 359 85
rect 359 67 375 85
rect 375 67 376 85
rect 463 95 465 113
rect 465 95 479 113
rect 479 95 481 113
rect 435 83 438 85
rect 438 83 452 85
rect 452 83 453 85
rect 560 84 578 102
rect 435 67 453 83
rect 532 56 550 74
<< metal2 >>
rect 84 526 96 758
rect 255 701 306 717
rect 532 715 544 758
rect 255 692 273 701
rect 532 698 550 715
rect 218 636 306 654
rect 324 636 406 654
rect 218 602 308 620
rect 192 574 227 592
rect 245 574 281 592
rect 299 574 431 592
rect 84 0 96 508
rect 127 347 139 548
rect 192 522 225 540
rect 243 522 297 540
rect 315 522 350 540
rect 368 522 430 540
rect 448 522 510 540
rect 217 494 324 512
rect 421 494 458 512
rect 324 475 342 494
rect 324 457 424 475
rect 538 361 550 698
rect 127 329 130 347
rect 127 177 139 329
rect 192 217 225 235
rect 243 217 359 235
rect 405 217 509 235
rect 270 189 413 207
rect 351 137 463 155
rect 244 95 305 113
rect 351 95 463 113
rect 376 67 435 85
rect 538 74 550 343
rect 560 102 572 758
rect 532 0 544 56
rect 560 0 572 84
<< labels >>
rlabel metal1 0 6 0 30 3 GND!
rlabel metal2 84 0 96 0 1 D
rlabel metal2 532 0 544 0 1 Q
rlabel metal2 560 0 572 0 1 nQ
rlabel metal1 588 263 588 273 7 nReset
rlabel metal1 588 288 588 298 7 Clock
rlabel metal1 588 307 588 317 7 Test
rlabel metal1 588 351 588 361 7 Q
rlabel metal1 588 370 588 380 7 ScanReturn
rlabel metal1 588 728 588 752 7 Vdd!
rlabel metal2 560 758 572 758 5 nQ
rlabel metal2 532 758 544 758 5 Q
rlabel metal1 0 263 0 273 3 nReset
rlabel metal1 0 288 0 298 3 Clock
rlabel metal1 0 307 0 317 3 Test
rlabel metal1 0 351 0 361 3 SDI
rlabel metal1 0 370 0 380 3 ScanReturn
rlabel metal1 0 728 0 752 3 Vdd!
rlabel metal2 84 758 96 758 5 D
rlabel metal1 588 6 588 30 7 GND!
<< end >>
