magic
tech c35b4
timestamp 1543772271
<< pimplant >>
rect 0 334 644 727
<< nimplant >>
rect 0 31 644 281
<< nwell >>
rect 0 334 644 752
<< polysilicon >>
rect 23 715 30 724
rect 23 593 30 659
rect 51 593 58 724
rect 79 715 86 724
rect 79 593 86 659
rect 107 593 114 724
rect 135 695 142 724
rect 135 593 142 679
rect 163 656 170 724
rect 163 593 170 640
rect 190 593 197 724
rect 247 624 254 727
rect 275 692 282 727
rect 303 692 310 727
rect 356 717 363 727
rect 356 701 362 717
rect 356 692 363 701
rect 389 692 396 727
rect 428 692 435 727
rect 481 692 488 727
rect 275 624 282 636
rect 303 571 310 636
rect 356 624 363 636
rect 247 540 254 568
rect 275 555 282 568
rect 303 564 335 571
rect 275 548 307 555
rect 300 540 307 548
rect 23 176 30 537
rect 51 219 58 537
rect 79 323 86 537
rect 107 364 114 537
rect 51 218 62 219
rect 51 201 62 202
rect 23 150 30 160
rect 51 150 58 201
rect 79 150 86 307
rect 107 150 114 348
rect 135 150 142 537
rect 163 150 170 537
rect 190 364 197 537
rect 196 348 197 364
rect 190 150 197 348
rect 247 298 254 484
rect 300 374 307 484
rect 275 367 307 374
rect 247 235 254 282
rect 275 279 282 367
rect 328 358 335 564
rect 356 555 363 568
rect 389 555 396 636
rect 428 624 435 636
rect 481 624 488 636
rect 428 560 435 568
rect 303 351 335 358
rect 344 548 363 555
rect 372 548 396 555
rect 425 553 435 560
rect 481 555 488 568
rect 514 567 521 727
rect 303 342 310 351
rect 303 303 310 326
rect 303 296 335 303
rect 275 247 282 263
rect 275 240 307 247
rect 300 235 307 240
rect 247 155 254 205
rect 300 200 307 205
rect 275 193 307 200
rect 275 155 282 193
rect 23 73 30 120
rect 23 34 30 43
rect 51 34 58 120
rect 79 73 86 120
rect 79 34 86 43
rect 107 34 114 120
rect 135 66 142 120
rect 163 92 170 120
rect 167 76 170 92
rect 135 34 142 50
rect 163 34 170 76
rect 190 34 197 120
rect 247 31 254 125
rect 275 113 282 125
rect 328 113 335 296
rect 344 166 351 548
rect 372 540 379 548
rect 425 540 432 553
rect 478 548 488 555
rect 505 549 514 556
rect 478 540 485 548
rect 505 540 512 549
rect 558 540 565 727
rect 372 358 379 484
rect 425 358 432 484
rect 478 475 485 484
rect 478 468 480 475
rect 485 358 492 457
rect 372 351 384 358
rect 425 351 442 358
rect 485 351 495 358
rect 377 235 384 351
rect 435 235 442 351
rect 488 235 495 351
rect 505 260 512 484
rect 558 475 565 484
rect 504 235 511 244
rect 557 235 564 459
rect 377 182 384 205
rect 377 175 422 182
rect 344 159 388 166
rect 381 155 388 159
rect 381 113 388 125
rect 415 85 422 175
rect 435 171 442 205
rect 488 180 495 205
rect 504 201 511 205
rect 504 194 546 201
rect 435 164 465 171
rect 504 164 518 171
rect 458 155 465 164
rect 511 155 518 164
rect 458 113 465 125
rect 511 113 518 125
rect 275 31 282 83
rect 328 31 335 83
rect 381 74 388 83
rect 381 31 388 58
rect 417 31 424 67
rect 458 31 465 83
rect 511 31 518 83
rect 539 74 546 194
rect 557 102 564 205
rect 539 31 546 56
rect 557 31 564 84
<< ndiffusion >>
rect 244 205 247 235
rect 254 205 257 235
rect 297 205 300 235
rect 307 205 310 235
rect 20 120 23 150
rect 30 120 51 150
rect 58 120 61 150
rect 75 120 79 150
rect 86 120 107 150
rect 114 120 118 150
rect 132 120 135 150
rect 142 120 145 150
rect 159 120 163 150
rect 170 120 190 150
rect 197 120 200 150
rect 244 125 247 155
rect 254 125 275 155
rect 282 125 285 155
rect 20 43 23 73
rect 30 43 33 73
rect 76 43 79 73
rect 86 43 89 73
rect 374 205 377 235
rect 384 205 392 235
rect 432 205 435 235
rect 442 205 445 235
rect 485 205 488 235
rect 495 205 504 235
rect 511 205 514 235
rect 554 205 557 235
rect 564 205 567 235
rect 378 125 381 155
rect 388 125 391 155
rect 272 83 275 113
rect 282 83 285 113
rect 325 83 328 113
rect 335 83 338 113
rect 378 83 381 113
rect 388 83 391 113
rect 508 125 511 155
rect 518 125 521 155
rect 455 83 458 113
rect 465 83 468 113
rect 508 83 511 113
rect 518 83 521 113
<< pdiffusion >>
rect 20 659 23 715
rect 30 659 33 715
rect 76 659 79 715
rect 86 659 89 715
rect 272 636 275 692
rect 282 636 285 692
rect 299 636 303 692
rect 310 636 313 692
rect 353 636 356 692
rect 363 636 366 692
rect 425 636 428 692
rect 435 636 438 692
rect 478 636 481 692
rect 488 636 491 692
rect 20 537 23 593
rect 30 537 34 593
rect 48 537 51 593
rect 58 537 61 593
rect 75 537 79 593
rect 86 537 89 593
rect 103 537 107 593
rect 114 537 118 593
rect 132 537 135 593
rect 142 537 146 593
rect 160 537 163 593
rect 170 537 173 593
rect 187 537 190 593
rect 197 537 201 593
rect 244 568 247 624
rect 254 568 257 624
rect 272 568 275 624
rect 282 568 285 624
rect 353 568 356 624
rect 363 568 366 624
rect 244 484 247 540
rect 254 484 257 540
rect 297 484 300 540
rect 307 484 310 540
rect 478 568 481 624
rect 488 568 491 624
rect 369 484 372 540
rect 379 484 382 540
rect 422 484 425 540
rect 432 484 435 540
rect 475 484 478 540
rect 485 484 488 540
rect 502 484 505 540
rect 512 484 515 540
rect 555 484 558 540
rect 565 484 568 540
<< ntransistor >>
rect 247 205 254 235
rect 300 205 307 235
rect 23 120 30 150
rect 51 120 58 150
rect 79 120 86 150
rect 107 120 114 150
rect 135 120 142 150
rect 163 120 170 150
rect 190 120 197 150
rect 247 125 254 155
rect 275 125 282 155
rect 23 43 30 73
rect 79 43 86 73
rect 377 205 384 235
rect 435 205 442 235
rect 488 205 495 235
rect 504 205 511 235
rect 557 205 564 235
rect 381 125 388 155
rect 275 83 282 113
rect 328 83 335 113
rect 381 83 388 113
rect 511 125 518 155
rect 458 83 465 113
rect 511 83 518 113
<< ptransistor >>
rect 23 659 30 715
rect 79 659 86 715
rect 275 636 282 692
rect 303 636 310 692
rect 356 636 363 692
rect 428 636 435 692
rect 481 636 488 692
rect 23 537 30 593
rect 51 537 58 593
rect 79 537 86 593
rect 107 537 114 593
rect 135 537 142 593
rect 163 537 170 593
rect 190 537 197 593
rect 247 568 254 624
rect 275 568 282 624
rect 356 568 363 624
rect 247 484 254 540
rect 300 484 307 540
rect 481 568 488 624
rect 372 484 379 540
rect 425 484 432 540
rect 478 484 485 540
rect 505 484 512 540
rect 558 484 565 540
<< polycontact >>
rect 126 679 142 695
rect 154 640 170 656
rect 362 701 378 717
rect 384 636 400 692
rect 107 348 123 364
rect 79 307 95 323
rect 51 202 67 218
rect 19 160 35 176
rect 180 348 196 364
rect 243 282 259 298
rect 428 568 444 624
rect 298 326 314 342
rect 271 263 287 279
rect 151 76 167 92
rect 131 50 147 66
rect 514 549 530 567
rect 480 457 496 475
rect 555 459 571 475
rect 504 244 520 260
rect 488 164 504 180
rect 449 125 465 155
rect 378 58 394 74
rect 415 67 431 85
rect 555 84 571 102
rect 530 56 546 74
<< ndiffcontact >>
rect 230 205 244 235
rect 257 205 271 235
rect 283 205 297 235
rect 310 205 324 235
rect 6 120 20 150
rect 61 120 75 150
rect 118 120 132 150
rect 145 120 159 150
rect 200 120 214 150
rect 230 125 244 155
rect 285 125 299 155
rect 6 43 20 73
rect 33 43 47 73
rect 62 43 76 73
rect 89 43 103 73
rect 360 205 374 235
rect 392 205 406 235
rect 418 205 432 235
rect 445 205 459 235
rect 471 205 485 235
rect 514 205 528 235
rect 540 205 554 235
rect 567 205 581 235
rect 364 125 378 155
rect 391 125 405 155
rect 258 83 272 113
rect 285 83 299 113
rect 311 83 325 113
rect 338 83 352 113
rect 364 83 378 113
rect 391 83 405 113
rect 494 125 508 155
rect 521 125 535 155
rect 441 83 455 113
rect 468 83 482 113
rect 494 83 508 113
rect 521 83 535 113
<< pdiffcontact >>
rect 6 659 20 715
rect 33 659 47 715
rect 62 659 76 715
rect 89 659 103 715
rect 258 636 272 692
rect 285 636 299 692
rect 313 636 327 692
rect 339 636 353 692
rect 366 636 380 692
rect 411 636 425 692
rect 438 636 452 692
rect 464 636 478 692
rect 491 636 505 692
rect 6 537 20 593
rect 34 537 48 593
rect 61 537 75 593
rect 89 537 103 593
rect 118 537 132 593
rect 146 537 160 593
rect 173 537 187 593
rect 201 537 215 593
rect 230 568 244 624
rect 257 568 272 624
rect 285 568 299 624
rect 339 568 353 624
rect 366 568 380 624
rect 230 484 244 540
rect 257 484 271 540
rect 283 484 297 540
rect 310 484 324 540
rect 464 568 478 624
rect 491 568 505 624
rect 355 484 369 540
rect 382 484 396 540
rect 408 484 422 540
rect 435 484 449 540
rect 461 484 475 540
rect 488 484 502 540
rect 515 484 529 540
rect 541 484 555 540
rect 568 484 582 540
<< psubstratetap >>
rect 6 10 638 24
<< nsubstratetap >>
rect 6 734 638 748
<< metal1 >>
rect 0 748 644 752
rect 0 734 6 748
rect 638 734 644 748
rect 0 728 644 734
rect 6 715 20 728
rect 62 715 76 728
rect 103 682 126 692
rect 35 650 45 659
rect 35 640 154 650
rect 36 621 185 631
rect 36 593 46 621
rect 63 602 130 612
rect 63 593 73 602
rect 120 593 130 602
rect 175 593 185 621
rect 201 593 215 728
rect 230 624 244 728
rect 285 692 299 728
rect 339 692 353 728
rect 380 701 425 717
rect 411 692 425 701
rect 380 636 384 692
rect 438 692 452 728
rect 491 692 505 728
rect 380 620 428 624
rect 382 602 428 620
rect 380 568 428 602
rect 444 568 464 624
rect 230 540 244 568
rect 435 549 514 559
rect 530 549 555 559
rect 435 540 449 549
rect 541 540 555 549
rect 8 528 18 537
rect 63 528 73 537
rect 8 518 73 528
rect 148 528 158 537
rect 203 528 213 537
rect 148 518 213 528
rect 310 475 324 484
rect 461 475 471 484
rect 515 475 529 484
rect 310 465 471 475
rect 515 459 555 475
rect 21 380 215 383
rect 0 373 644 380
rect 0 370 31 373
rect 205 370 644 373
rect 0 351 107 361
rect 196 351 588 361
rect 606 351 644 361
rect 171 329 298 339
rect 0 307 79 317
rect 95 307 644 317
rect 0 288 243 298
rect 259 288 644 298
rect 0 263 271 273
rect 456 273 554 279
rect 287 269 644 273
rect 287 263 466 269
rect 544 263 644 269
rect 257 244 374 254
rect 520 244 554 254
rect 257 235 271 244
rect 360 235 374 244
rect 540 235 554 244
rect 63 182 194 192
rect 63 150 73 182
rect 118 159 190 173
rect 118 150 132 159
rect 8 111 18 120
rect 147 111 157 120
rect 8 101 157 111
rect 35 82 151 92
rect 35 73 45 82
rect 103 53 131 63
rect 6 30 20 43
rect 62 30 76 43
rect 176 30 190 159
rect 202 150 212 182
rect 230 155 244 205
rect 392 174 406 205
rect 514 196 528 205
rect 514 186 571 196
rect 392 164 488 174
rect 299 125 364 155
rect 465 125 494 155
rect 230 113 244 125
rect 230 83 258 113
rect 230 30 244 83
rect 311 49 325 83
rect 338 74 352 83
rect 338 58 378 74
rect 441 49 455 83
rect 311 39 455 49
rect 555 102 571 186
rect 468 30 482 83
rect 571 84 616 102
rect 546 56 588 74
rect 0 24 644 30
rect 0 10 6 24
rect 638 10 644 24
rect 0 6 644 10
<< m2contact >>
rect 87 537 89 555
rect 89 537 103 555
rect 103 537 105 555
rect 362 717 380 719
rect 362 701 378 717
rect 378 701 380 717
rect 256 636 258 654
rect 258 636 272 654
rect 272 636 274 654
rect 311 674 313 692
rect 313 674 327 692
rect 327 674 329 692
rect 362 636 366 654
rect 366 636 380 654
rect 462 636 464 654
rect 464 636 478 654
rect 478 636 480 654
rect 256 602 257 620
rect 257 602 272 620
rect 272 602 274 620
rect 230 574 244 592
rect 244 574 248 592
rect 364 602 366 620
rect 366 602 380 620
rect 380 602 382 620
rect 283 574 285 592
rect 285 574 299 592
rect 299 574 301 592
rect 337 574 339 592
rect 339 574 353 592
rect 353 574 355 592
rect 487 574 491 592
rect 491 574 505 592
rect 230 522 244 540
rect 244 522 248 540
rect 281 522 283 540
rect 283 522 297 540
rect 297 522 299 540
rect 255 494 257 512
rect 257 494 271 512
rect 271 494 273 512
rect 353 522 355 540
rect 355 522 369 540
rect 369 522 371 540
rect 406 522 408 540
rect 408 522 422 540
rect 422 522 424 540
rect 380 494 382 512
rect 382 494 396 512
rect 396 494 398 512
rect 486 522 488 540
rect 488 522 502 540
rect 502 522 504 540
rect 459 494 461 512
rect 461 494 475 512
rect 475 494 477 512
rect 514 494 515 512
rect 515 494 529 512
rect 529 494 532 512
rect 566 522 568 540
rect 568 522 582 540
rect 582 522 584 540
rect 480 457 496 475
rect 496 457 498 475
rect 153 329 171 347
rect 588 343 606 361
rect 50 218 68 219
rect 50 202 51 218
rect 51 202 67 218
rect 67 202 68 218
rect 50 201 68 202
rect 230 217 244 235
rect 244 217 248 235
rect 281 217 283 235
rect 283 217 297 235
rect 297 217 299 235
rect 308 205 310 207
rect 310 205 324 207
rect 324 205 326 207
rect 415 217 418 235
rect 418 217 432 235
rect 432 217 433 235
rect 443 217 445 235
rect 445 217 459 235
rect 459 217 461 235
rect 469 205 471 207
rect 471 205 485 207
rect 485 205 487 207
rect 194 182 212 200
rect 18 176 36 177
rect 18 160 19 176
rect 19 160 35 176
rect 35 160 36 176
rect 18 159 36 160
rect 308 189 326 205
rect 469 189 487 205
rect 565 217 567 235
rect 567 217 581 235
rect 581 217 583 235
rect 389 137 391 155
rect 391 137 405 155
rect 405 137 407 155
rect 519 137 521 155
rect 521 137 535 155
rect 535 137 537 155
rect 282 95 285 113
rect 285 95 299 113
rect 299 95 300 113
rect 361 95 364 113
rect 364 95 378 113
rect 378 95 379 113
rect 389 95 391 113
rect 391 95 405 113
rect 405 95 407 113
rect 414 67 415 85
rect 415 67 431 85
rect 431 67 432 85
rect 519 95 521 113
rect 521 95 535 113
rect 535 95 537 113
rect 491 83 494 85
rect 494 83 508 85
rect 508 83 509 85
rect 616 84 634 102
rect 491 67 509 83
rect 588 56 606 74
<< metal2 >>
rect 28 177 40 758
rect 56 219 68 758
rect 311 701 362 717
rect 588 715 600 758
rect 311 692 329 701
rect 588 698 606 715
rect 274 636 362 654
rect 380 636 462 654
rect 274 602 364 620
rect 248 574 283 592
rect 301 574 337 592
rect 355 574 487 592
rect 90 344 102 537
rect 248 522 281 540
rect 299 522 353 540
rect 371 522 406 540
rect 424 522 486 540
rect 504 522 566 540
rect 273 494 380 512
rect 477 494 514 512
rect 380 475 398 494
rect 380 457 480 475
rect 594 361 606 698
rect 90 332 153 344
rect 171 330 209 342
rect 36 159 40 177
rect 28 0 40 159
rect 56 0 68 201
rect 197 200 209 330
rect 248 217 281 235
rect 299 217 415 235
rect 461 217 565 235
rect 326 189 469 207
rect 407 137 519 155
rect 300 95 361 113
rect 407 95 519 113
rect 432 67 491 85
rect 594 74 606 343
rect 616 102 628 758
rect 588 0 600 56
rect 616 0 628 84
<< labels >>
rlabel metal1 0 728 0 752 3 Vdd!
rlabel metal2 28 758 40 758 5 Load
rlabel metal2 56 758 68 758 5 D
rlabel metal2 588 758 600 758 5 Q
rlabel metal2 616 758 628 758 5 nQ
rlabel metal1 644 728 644 752 7 Vdd!
rlabel metal1 644 263 644 273 7 nReset
rlabel metal1 644 288 644 298 7 Clock
rlabel metal1 644 307 644 317 7 Test
rlabel metal1 644 351 644 361 7 Q
rlabel metal1 644 370 644 380 7 ScanReturn
rlabel metal1 644 6 644 30 7 GND!
rlabel metal2 588 0 600 0 1 Q
rlabel metal2 616 0 628 0 1 nQ
rlabel metal2 56 0 68 0 1 D
rlabel metal2 28 0 40 0 1 Load
rlabel metal1 0 6 0 30 3 GND!
rlabel metal1 0 263 0 273 3 nReset
rlabel metal1 0 288 0 298 3 Clock
rlabel metal1 0 307 0 317 3 Test
rlabel metal1 0 351 0 361 3 SDI
rlabel metal1 0 370 0 380 3 ScanReturn
<< end >>
