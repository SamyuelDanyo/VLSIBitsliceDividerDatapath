magic
tech c35b4
timestamp 1543772418
<< pimplant >>
rect 0 334 140 727
<< nimplant >>
rect 0 31 140 281
<< nwell >>
rect 0 334 140 752
<< polysilicon >>
rect 23 719 30 727
rect 50 719 57 727
rect 77 719 84 727
rect 23 96 30 663
rect 50 96 57 663
rect 77 96 84 663
rect 23 69 30 78
rect 50 69 57 78
rect 77 69 84 78
rect 23 31 30 39
rect 50 31 57 39
rect 77 31 84 39
<< ndiffusion >>
rect 20 39 23 69
rect 30 39 50 69
rect 57 39 77 69
rect 84 39 87 69
<< pdiffusion >>
rect 20 663 23 719
rect 30 663 33 719
rect 47 663 50 719
rect 57 663 60 719
rect 74 663 77 719
rect 84 663 87 719
<< ntransistor >>
rect 23 39 30 69
rect 50 39 57 69
rect 77 39 84 69
<< ptransistor >>
rect 23 663 30 719
rect 50 663 57 719
rect 77 663 84 719
<< polycontact >>
rect 23 78 39 96
rect 50 78 68 96
rect 77 78 95 96
<< ndiffcontact >>
rect 6 39 20 69
rect 87 39 101 69
<< pdiffcontact >>
rect 6 663 20 719
rect 33 663 47 719
rect 60 663 74 719
rect 87 663 101 719
<< psubstratetap >>
rect 6 10 134 24
<< nsubstratetap >>
rect 6 734 134 748
<< metal1 >>
rect 0 748 140 752
rect 0 734 6 748
rect 134 734 140 748
rect 0 728 140 734
rect 6 719 20 728
rect 60 719 74 728
rect 101 663 106 719
rect 33 654 47 663
rect 87 654 101 663
rect 33 644 101 654
rect 0 370 140 380
rect 0 351 140 361
rect 0 307 140 317
rect 0 288 140 298
rect 0 263 140 273
rect 101 39 106 69
rect 6 30 20 39
rect 0 24 140 30
rect 0 10 6 24
rect 134 10 140 24
rect 0 6 140 10
<< m2contact >>
rect 106 663 124 719
rect 22 78 23 96
rect 23 78 39 96
rect 39 78 40 96
rect 50 78 68 96
rect 78 78 95 96
rect 95 78 96 96
rect 106 39 124 69
<< metal2 >>
rect 28 96 40 758
rect 56 96 68 758
rect 84 96 96 758
rect 112 719 124 758
rect 28 0 40 78
rect 56 0 68 78
rect 84 0 96 78
rect 112 69 124 663
rect 112 0 124 39
<< labels >>
rlabel metal2 28 0 40 0 1 A
rlabel metal2 56 0 68 0 1 B
rlabel metal2 84 0 96 0 1 C
rlabel metal2 112 0 124 0 1 Y
rlabel metal1 0 6 0 30 3 GND!
rlabel metal1 140 6 140 30 7 GND!
rlabel metal2 112 758 124 758 5 Y
rlabel metal2 84 758 96 758 5 C
rlabel metal2 56 758 68 758 5 B
rlabel metal2 28 758 40 758 5 A
rlabel metal1 0 728 0 752 3 Vdd!
rlabel metal1 140 728 140 752 7 Vdd!
rlabel metal1 0 263 0 273 3 nReset
rlabel metal1 0 307 0 317 3 Test
rlabel metal1 0 288 0 298 3 Clock
rlabel metal1 0 370 0 380 3 ScanReturn
rlabel metal1 0 351 0 361 3 Scan
rlabel metal1 140 263 140 273 7 nReset
rlabel metal1 140 288 140 298 7 Clock
rlabel metal1 140 307 140 317 7 Test
rlabel metal1 140 351 140 361 7 Scan
rlabel metal1 140 370 140 380 7 ScanReturn
<< end >>
