magic
tech c35b4
timestamp 1547137389
<< metal1 >>
rect 0 84 305 94
rect 0 56 5386 66
rect 5376 38 5386 56
rect 0 28 5358 38
rect 5376 28 5554 38
rect 5348 15 5358 28
rect 5544 15 5554 28
rect 392 -830 402 -815
rect 252 -840 402 -830
rect 252 -914 262 -840
rect 7112 -830 7122 -815
rect 435 -840 7122 -830
rect 7756 -830 7766 -815
rect 7155 -840 7766 -830
rect 8176 -830 8186 -815
rect 7799 -840 8186 -830
rect 8288 -830 8298 -815
rect 8247 -840 8298 -830
rect 280 -868 5569 -858
rect 280 -909 290 -868
rect 5587 -868 8061 -858
rect 8079 -868 8257 -858
rect 392 -896 5065 -886
rect 392 -909 402 -896
rect 5111 -896 6073 -886
rect 6119 -896 6941 -886
rect 6987 -896 7697 -886
rect 7715 -896 8145 -886
rect 8191 -896 8229 -886
rect 224 -924 262 -914
rect 224 -1189 234 -924
rect 463 -924 5849 -914
rect 5895 -924 6409 -914
rect 6455 -924 7473 -914
rect 7491 -924 7837 -914
rect 7911 -924 8201 -914
rect 252 -952 5961 -942
rect 252 -1189 262 -952
rect 6007 -952 6857 -942
rect 6903 -952 8089 -942
rect 8120 -952 8173 -942
rect 476 -980 7949 -970
rect 280 -1189 290 -983
rect 308 -1222 318 -983
rect 336 -1217 346 -983
rect 168 -1232 318 -1222
rect 168 -1278 178 -1232
rect 364 -1250 374 -983
rect 392 -1245 402 -983
rect 420 -1245 430 -983
rect 448 -1245 458 -983
rect 196 -1260 374 -1250
rect 196 -1273 206 -1260
rect 140 -1288 178 -1278
rect 140 -1357 150 -1288
rect 476 -1278 486 -980
rect 8023 -980 8033 -970
rect 8120 -970 8130 -952
rect 8064 -980 8130 -970
rect 1443 -1008 2013 -998
rect 2059 -1008 5485 -998
rect 5531 -1008 5681 -998
rect 5699 -1008 5821 -998
rect 5839 -1008 6045 -998
rect 6063 -1008 6269 -998
rect 6287 -1008 6493 -998
rect 6511 -1008 7277 -998
rect 7323 -1008 7865 -998
rect 8064 -998 8074 -980
rect 7939 -1008 8074 -998
rect 1891 -1036 4701 -1026
rect 4719 -1036 4953 -1026
rect 4971 -1036 7613 -1026
rect 7687 -1036 7725 -1026
rect 7771 -1036 8005 -1026
rect 1919 -1064 5457 -1054
rect 5503 -1064 6185 -1054
rect 6231 -1064 6241 -1054
rect 6259 -1064 6353 -1054
rect 6371 -1064 7025 -1054
rect 7071 -1064 7977 -1054
rect 1975 -1092 4729 -1082
rect 4775 -1092 5261 -1082
rect 5307 -1092 6633 -1082
rect 6679 -1092 7389 -1082
rect 7435 -1092 7809 -1082
rect 7840 -1092 7893 -1082
rect 2003 -1120 2041 -1110
rect 2143 -1120 4617 -1110
rect 7840 -1110 7850 -1092
rect 4663 -1120 7850 -1110
rect 2591 -1148 4897 -1138
rect 4915 -1148 5401 -1138
rect 5419 -1148 7333 -1138
rect 7351 -1148 7557 -1138
rect 7575 -1148 7781 -1138
rect 2619 -1176 5709 -1166
rect 5783 -1176 7753 -1166
rect 2731 -1204 4841 -1194
rect 4887 -1204 6745 -1194
rect 6791 -1204 7165 -1194
rect 7183 -1204 7501 -1194
rect 7547 -1204 7641 -1194
rect 3179 -1232 6717 -1222
rect 6735 -1232 7585 -1222
rect 7672 -1222 7682 -1207
rect 7616 -1232 7682 -1222
rect 3207 -1260 7361 -1250
rect 7407 -1260 7445 -1250
rect 7616 -1250 7626 -1232
rect 7463 -1260 7626 -1250
rect 323 -1288 486 -1278
rect 3319 -1288 3889 -1278
rect 3935 -1288 6521 -1278
rect 6567 -1288 6997 -1278
rect 7015 -1288 7529 -1278
rect 168 -1316 333 -1306
rect 168 -1357 178 -1316
rect 379 -1316 417 -1306
rect 3767 -1316 6381 -1306
rect 6399 -1316 6605 -1306
rect 6623 -1316 7417 -1306
rect 448 -1334 458 -1319
rect 336 -1344 458 -1334
rect 196 -1357 206 -1347
rect 224 -1357 234 -1347
rect 252 -1357 262 -1347
rect 280 -1357 290 -1347
rect 308 -1357 318 -1347
rect 336 -1357 346 -1344
rect 3795 -1344 6829 -1334
rect 6847 -1344 7389 -1334
rect 3851 -1372 5625 -1362
rect 5671 -1372 6157 -1362
rect 6175 -1372 7193 -1362
rect 7267 -1372 7305 -1362
rect 3879 -1400 3917 -1390
rect 4019 -1400 5149 -1390
rect 5195 -1400 6297 -1390
rect 6343 -1400 6913 -1390
rect 6931 -1400 7053 -1390
rect 7099 -1400 7137 -1390
rect 4467 -1428 6969 -1418
rect 4495 -1456 5233 -1446
rect 5251 -1456 5933 -1446
rect 5951 -1456 6437 -1446
rect 6483 -1456 6549 -1446
rect 6595 -1456 6661 -1446
rect 6707 -1456 6773 -1446
rect 6819 -1456 6885 -1446
rect 4551 -1484 5737 -1474
rect 5811 -1484 6325 -1474
rect 4579 -1512 5877 -1502
rect 5923 -1512 5989 -1502
rect 6035 -1512 6101 -1502
rect 6147 -1512 6213 -1502
rect 4607 -1540 4645 -1530
rect 4691 -1540 4757 -1530
rect 4803 -1540 4981 -1530
rect 5012 -1540 5429 -1530
rect 4831 -1568 4869 -1558
rect 5012 -1558 5022 -1540
rect 5447 -1540 5513 -1530
rect 5559 -1540 5765 -1530
rect 4943 -1568 5022 -1558
rect 5055 -1568 5093 -1558
rect 5139 -1568 5177 -1558
rect 5223 -1568 5289 -1558
rect 5335 -1568 5485 -1558
rect 5615 -1568 5653 -1558
<< m2contact >>
rect 305 81 323 99
rect 5345 -3 5363 15
rect 5541 -3 5559 15
rect 389 -815 407 -797
rect 7109 -815 7127 -797
rect 7753 -815 7771 -797
rect 8173 -815 8191 -797
rect 8285 -815 8303 -797
rect 417 -843 435 -825
rect 7137 -843 7155 -825
rect 7781 -843 7799 -825
rect 8201 -843 8219 -825
rect 8229 -843 8247 -825
rect 5569 -871 5587 -853
rect 8061 -871 8079 -853
rect 8257 -871 8275 -853
rect 5065 -899 5083 -881
rect 5093 -899 5111 -881
rect 6073 -899 6091 -881
rect 6101 -899 6119 -881
rect 6941 -899 6959 -881
rect 6969 -899 6987 -881
rect 7697 -899 7715 -881
rect 8145 -899 8163 -881
rect 8173 -899 8191 -881
rect 8229 -899 8247 -881
rect 277 -927 295 -909
rect 389 -927 407 -909
rect 445 -927 463 -909
rect 5849 -927 5867 -909
rect 5877 -927 5895 -909
rect 6409 -927 6427 -909
rect 6437 -927 6455 -909
rect 7473 -927 7491 -909
rect 7837 -927 7855 -909
rect 7893 -927 7911 -909
rect 8201 -927 8219 -909
rect 5961 -955 5979 -937
rect 5989 -955 6007 -937
rect 6857 -955 6875 -937
rect 6885 -955 6903 -937
rect 8089 -955 8107 -937
rect 277 -983 295 -965
rect 305 -983 323 -965
rect 333 -983 351 -965
rect 361 -983 379 -965
rect 389 -983 407 -965
rect 417 -983 435 -965
rect 445 -983 463 -965
rect 221 -1207 239 -1189
rect 249 -1207 267 -1189
rect 277 -1207 295 -1189
rect 333 -1235 351 -1217
rect 389 -1263 407 -1245
rect 417 -1263 435 -1245
rect 445 -1263 463 -1245
rect 193 -1291 211 -1273
rect 305 -1291 323 -1273
rect 7949 -983 7967 -965
rect 8005 -983 8023 -965
rect 8033 -983 8051 -965
rect 8173 -955 8191 -937
rect 1425 -1011 1443 -993
rect 2013 -1011 2031 -993
rect 2041 -1011 2059 -993
rect 5485 -1011 5503 -993
rect 5513 -1011 5531 -993
rect 5681 -1011 5699 -993
rect 5821 -1011 5839 -993
rect 6045 -1011 6063 -993
rect 6269 -1011 6287 -993
rect 6493 -1011 6511 -993
rect 7277 -1011 7295 -993
rect 7305 -1011 7323 -993
rect 7865 -1011 7883 -993
rect 7921 -1011 7939 -993
rect 1873 -1039 1891 -1021
rect 4701 -1039 4719 -1021
rect 4953 -1039 4971 -1021
rect 7613 -1039 7631 -1021
rect 7669 -1039 7687 -1021
rect 7725 -1039 7743 -1021
rect 7753 -1039 7771 -1021
rect 8005 -1039 8023 -1021
rect 1901 -1067 1919 -1049
rect 5457 -1067 5475 -1049
rect 5485 -1067 5503 -1049
rect 6185 -1067 6203 -1049
rect 6213 -1067 6231 -1049
rect 6241 -1067 6259 -1049
rect 6353 -1067 6371 -1049
rect 7025 -1067 7043 -1049
rect 7053 -1067 7071 -1049
rect 7977 -1067 7995 -1049
rect 1957 -1095 1975 -1077
rect 4729 -1095 4747 -1077
rect 4757 -1095 4775 -1077
rect 5261 -1095 5279 -1077
rect 5289 -1095 5307 -1077
rect 6633 -1095 6651 -1077
rect 6661 -1095 6679 -1077
rect 7389 -1095 7407 -1077
rect 7417 -1095 7435 -1077
rect 7809 -1095 7827 -1077
rect 1985 -1123 2003 -1105
rect 2041 -1123 2059 -1105
rect 2125 -1123 2143 -1105
rect 4617 -1123 4635 -1105
rect 4645 -1123 4663 -1105
rect 7893 -1095 7911 -1077
rect 2573 -1151 2591 -1133
rect 4897 -1151 4915 -1133
rect 5401 -1151 5419 -1133
rect 7333 -1151 7351 -1133
rect 7557 -1151 7575 -1133
rect 7781 -1151 7799 -1133
rect 2601 -1179 2619 -1161
rect 5709 -1179 5727 -1161
rect 5765 -1179 5783 -1161
rect 7753 -1179 7771 -1161
rect 2713 -1207 2731 -1189
rect 4841 -1207 4859 -1189
rect 4869 -1207 4887 -1189
rect 6745 -1207 6763 -1189
rect 6773 -1207 6791 -1189
rect 7165 -1207 7183 -1189
rect 7501 -1207 7519 -1189
rect 7529 -1207 7547 -1189
rect 7641 -1207 7659 -1189
rect 7669 -1207 7687 -1189
rect 3161 -1235 3179 -1217
rect 6717 -1235 6735 -1217
rect 7585 -1235 7603 -1217
rect 3189 -1263 3207 -1245
rect 7361 -1263 7379 -1245
rect 7389 -1263 7407 -1245
rect 7445 -1263 7463 -1245
rect 3301 -1291 3319 -1273
rect 3889 -1291 3907 -1273
rect 3917 -1291 3935 -1273
rect 6521 -1291 6539 -1273
rect 6549 -1291 6567 -1273
rect 6997 -1291 7015 -1273
rect 7529 -1291 7547 -1273
rect 333 -1319 351 -1301
rect 361 -1319 379 -1301
rect 417 -1319 435 -1301
rect 445 -1319 463 -1301
rect 3749 -1319 3767 -1301
rect 6381 -1319 6399 -1301
rect 6605 -1319 6623 -1301
rect 7417 -1319 7435 -1301
rect 193 -1347 211 -1329
rect 221 -1347 239 -1329
rect 249 -1347 267 -1329
rect 277 -1347 295 -1329
rect 305 -1347 323 -1329
rect 3777 -1347 3795 -1329
rect 6829 -1347 6847 -1329
rect 7389 -1347 7407 -1329
rect 137 -1375 155 -1357
rect 165 -1375 183 -1357
rect 193 -1375 211 -1357
rect 221 -1375 239 -1357
rect 249 -1375 267 -1357
rect 277 -1375 295 -1357
rect 305 -1375 323 -1357
rect 333 -1375 351 -1357
rect 3833 -1375 3851 -1357
rect 5625 -1375 5643 -1357
rect 5653 -1375 5671 -1357
rect 6157 -1375 6175 -1357
rect 7193 -1375 7211 -1357
rect 7249 -1375 7267 -1357
rect 7305 -1375 7323 -1357
rect 3861 -1403 3879 -1385
rect 3917 -1403 3935 -1385
rect 4001 -1403 4019 -1385
rect 5149 -1403 5167 -1385
rect 5177 -1403 5195 -1385
rect 6297 -1403 6315 -1385
rect 6325 -1403 6343 -1385
rect 6913 -1403 6931 -1385
rect 7053 -1403 7071 -1385
rect 7081 -1403 7099 -1385
rect 7137 -1403 7155 -1385
rect 4449 -1431 4467 -1413
rect 6969 -1431 6987 -1413
rect 4477 -1459 4495 -1441
rect 5233 -1459 5251 -1441
rect 5933 -1459 5951 -1441
rect 6437 -1459 6455 -1441
rect 6465 -1459 6483 -1441
rect 6549 -1459 6567 -1441
rect 6577 -1459 6595 -1441
rect 6661 -1459 6679 -1441
rect 6689 -1459 6707 -1441
rect 6773 -1459 6791 -1441
rect 6801 -1459 6819 -1441
rect 6885 -1459 6903 -1441
rect 4533 -1487 4551 -1469
rect 5737 -1487 5755 -1469
rect 5793 -1487 5811 -1469
rect 6325 -1487 6343 -1469
rect 4561 -1515 4579 -1497
rect 5877 -1515 5895 -1497
rect 5905 -1515 5923 -1497
rect 5989 -1515 6007 -1497
rect 6017 -1515 6035 -1497
rect 6101 -1515 6119 -1497
rect 6129 -1515 6147 -1497
rect 6213 -1515 6231 -1497
rect 4589 -1543 4607 -1525
rect 4645 -1543 4663 -1525
rect 4673 -1543 4691 -1525
rect 4757 -1543 4775 -1525
rect 4785 -1543 4803 -1525
rect 4981 -1543 4999 -1525
rect 4813 -1571 4831 -1553
rect 4869 -1571 4887 -1553
rect 4925 -1571 4943 -1553
rect 5429 -1543 5447 -1525
rect 5513 -1543 5531 -1525
rect 5541 -1543 5559 -1525
rect 5765 -1543 5783 -1525
rect 5037 -1571 5055 -1553
rect 5093 -1571 5111 -1553
rect 5121 -1571 5139 -1553
rect 5177 -1571 5195 -1553
rect 5205 -1571 5223 -1553
rect 5289 -1571 5307 -1553
rect 5317 -1571 5335 -1553
rect 5485 -1571 5503 -1553
rect 5597 -1571 5615 -1553
rect 5653 -1571 5671 -1553
<< metal2 >>
rect 308 -28 320 81
rect 5348 -28 5360 -3
rect 5544 -28 5556 -3
rect 280 -965 292 -927
rect 308 -965 320 -786
rect 336 -965 348 -786
rect 364 -965 376 -786
rect 392 -797 404 -786
rect 392 -965 404 -927
rect 420 -965 432 -843
rect 448 -965 460 -927
rect 1428 -993 1440 -786
rect 1876 -1021 1888 -786
rect 1904 -1049 1916 -786
rect 1960 -1077 1972 -786
rect 1988 -1105 2000 -786
rect 2016 -993 2028 -786
rect 2044 -1105 2056 -1011
rect 2128 -1105 2140 -786
rect 2576 -1133 2588 -786
rect 2604 -1161 2616 -786
rect 2716 -1189 2728 -786
rect 196 -1329 208 -1291
rect 224 -1329 236 -1207
rect 252 -1329 264 -1207
rect 280 -1329 292 -1207
rect 3164 -1217 3176 -786
rect 308 -1329 320 -1291
rect 336 -1301 348 -1235
rect 3192 -1245 3204 -786
rect 140 -1388 152 -1375
rect 168 -1388 180 -1375
rect 196 -1388 208 -1375
rect 224 -1388 236 -1375
rect 252 -1388 264 -1375
rect 280 -1388 292 -1375
rect 308 -1388 320 -1375
rect 336 -1388 348 -1375
rect 364 -1388 376 -1319
rect 392 -1388 404 -1263
rect 420 -1301 432 -1263
rect 448 -1301 460 -1263
rect 3304 -1273 3316 -786
rect 3752 -1301 3764 -786
rect 3780 -1329 3792 -786
rect 3836 -1357 3848 -786
rect 3864 -1385 3876 -786
rect 3892 -1273 3904 -786
rect 3920 -1385 3932 -1291
rect 4004 -1385 4016 -786
rect 4452 -1413 4464 -786
rect 4480 -1441 4492 -786
rect 4536 -1469 4548 -786
rect 4564 -1497 4576 -786
rect 4592 -1525 4604 -786
rect 4620 -1105 4632 -786
rect 4648 -1525 4660 -1123
rect 4676 -1525 4688 -786
rect 4704 -1021 4716 -786
rect 4732 -1077 4744 -786
rect 4760 -1525 4772 -1095
rect 4788 -1525 4800 -786
rect 4816 -1553 4828 -786
rect 4844 -1189 4856 -786
rect 4900 -1133 4912 -786
rect 4872 -1553 4884 -1207
rect 4928 -1553 4940 -786
rect 4956 -1021 4968 -786
rect 4984 -1525 4996 -786
rect 5040 -1553 5052 -786
rect 5068 -881 5080 -786
rect 5096 -1553 5108 -899
rect 5124 -1553 5136 -786
rect 5152 -1385 5164 -786
rect 5180 -1553 5192 -1403
rect 5208 -1553 5220 -786
rect 5236 -1441 5248 -786
rect 5264 -1077 5276 -786
rect 5292 -1553 5304 -1095
rect 5320 -1553 5332 -786
rect 5404 -1133 5416 -786
rect 5432 -1525 5444 -786
rect 5460 -1049 5472 -786
rect 5488 -993 5500 -786
rect 5488 -1553 5500 -1067
rect 5516 -1525 5528 -1011
rect 5544 -1525 5556 -786
rect 5572 -853 5584 -786
rect 5600 -1553 5612 -786
rect 5628 -1357 5640 -786
rect 5684 -993 5696 -786
rect 5712 -1161 5724 -786
rect 5656 -1553 5668 -1375
rect 5740 -1469 5752 -786
rect 5768 -1525 5780 -1179
rect 5796 -1469 5808 -786
rect 5824 -993 5836 -786
rect 5852 -909 5864 -786
rect 5880 -1497 5892 -927
rect 5908 -1497 5920 -786
rect 5936 -1441 5948 -786
rect 5964 -937 5976 -786
rect 5992 -1497 6004 -955
rect 6020 -1497 6032 -786
rect 6048 -993 6060 -786
rect 6076 -881 6088 -786
rect 6104 -1497 6116 -899
rect 6132 -1497 6144 -786
rect 6160 -1357 6172 -786
rect 6188 -1049 6200 -786
rect 6244 -1049 6256 -786
rect 6272 -993 6284 -786
rect 6216 -1497 6228 -1067
rect 6300 -1385 6312 -786
rect 6356 -1049 6368 -786
rect 6384 -1301 6396 -786
rect 6412 -909 6424 -786
rect 6328 -1469 6340 -1403
rect 6440 -1441 6452 -927
rect 6468 -1441 6480 -786
rect 6496 -993 6508 -786
rect 6524 -1273 6536 -786
rect 6552 -1441 6564 -1291
rect 6580 -1441 6592 -786
rect 6608 -1301 6620 -786
rect 6636 -1077 6648 -786
rect 6664 -1441 6676 -1095
rect 6692 -1441 6704 -786
rect 6720 -1217 6732 -786
rect 6748 -1189 6760 -786
rect 6776 -1441 6788 -1207
rect 6804 -1441 6816 -786
rect 6832 -1329 6844 -786
rect 6860 -937 6872 -786
rect 6888 -1441 6900 -955
rect 6916 -1385 6928 -786
rect 6944 -881 6956 -786
rect 6972 -1413 6984 -899
rect 7000 -1273 7012 -786
rect 7028 -1049 7040 -786
rect 7056 -1385 7068 -1067
rect 7084 -1385 7096 -786
rect 7112 -797 7124 -786
rect 7140 -1385 7152 -843
rect 7168 -1189 7180 -786
rect 7196 -1357 7208 -786
rect 7252 -1357 7264 -786
rect 7280 -993 7292 -786
rect 7308 -1357 7320 -1011
rect 7336 -1133 7348 -786
rect 7364 -1245 7376 -786
rect 7392 -1077 7404 -786
rect 7392 -1329 7404 -1263
rect 7420 -1301 7432 -1095
rect 7448 -1245 7460 -786
rect 7476 -909 7488 -786
rect 7504 -1189 7516 -786
rect 7560 -1133 7572 -786
rect 7532 -1273 7544 -1207
rect 7588 -1217 7600 -786
rect 7616 -1021 7628 -786
rect 7644 -1189 7656 -786
rect 7700 -881 7712 -786
rect 7728 -1021 7740 -786
rect 7756 -797 7768 -786
rect 7672 -1189 7684 -1039
rect 7756 -1161 7768 -1039
rect 7784 -1133 7796 -843
rect 7812 -1077 7824 -786
rect 7840 -909 7852 -786
rect 7868 -993 7880 -786
rect 7896 -1077 7908 -927
rect 7924 -993 7936 -786
rect 7952 -965 7964 -786
rect 7980 -1049 7992 -786
rect 8036 -965 8048 -786
rect 8064 -853 8076 -786
rect 8092 -937 8104 -786
rect 8148 -881 8160 -786
rect 8176 -797 8188 -786
rect 8204 -825 8216 -786
rect 8176 -937 8188 -899
rect 8204 -909 8216 -843
rect 8232 -881 8244 -843
rect 8260 -853 8272 -786
rect 8288 -797 8300 -786
rect 8008 -1021 8020 -983
use leftbuf  leftbuf_0
timestamp 1544089383
transform 1 0 28 0 1 -786
box 0 0 1316 758
use scandtype  cnt_reg_1
timestamp 1543772215
transform 1 0 1344 0 1 -786
box 0 0 588 758
use nand2  g602
timestamp 1543772396
transform 1 0 1932 0 1 -786
box 0 0 112 758
use scandtype  cnt_reg_0
timestamp 1543772215
transform 1 0 2044 0 1 -786
box 0 0 588 758
use scandtype  cnt_reg_2
timestamp 1543772215
transform 1 0 2632 0 1 -786
box 0 0 588 758
use scandtype  state_reg_0
timestamp 1543772215
transform 1 0 3220 0 1 -786
box 0 0 588 758
use nand2  g607
timestamp 1543772396
transform 1 0 3808 0 1 -786
box 0 0 112 758
use scandtype  state_reg_1
timestamp 1543772215
transform 1 0 3920 0 1 -786
box 0 0 588 758
use nand3  g603
timestamp 1543772418
transform 1 0 4508 0 1 -786
box 0 0 140 758
use nand2  g605
timestamp 1543772396
transform 1 0 4648 0 1 -786
box 0 0 112 758
use nand2  g615
timestamp 1543772396
transform 1 0 4760 0 1 -786
box 0 0 112 758
use nand3  g620
timestamp 1543772418
transform 1 0 4872 0 1 -786
box 0 0 140 758
use inv  g619
timestamp 1543772090
transform 1 0 5012 0 1 -786
box 0 0 84 758
use inv  g609
timestamp 1543772090
transform 1 0 5096 0 1 -786
box 0 0 84 758
use nand2  g614
timestamp 1543772396
transform 1 0 5180 0 1 -786
box 0 0 112 758
use inv  g610
timestamp 1543772090
transform 1 0 5292 0 1 -786
box 0 0 84 758
use nand3  g626
timestamp 1543772418
transform 1 0 5376 0 1 -786
box 0 0 140 758
use nand3  g618
timestamp 1543772418
transform 1 0 5516 0 1 -786
box 0 0 140 758
use nand2  g621
timestamp 1543772396
transform 1 0 5656 0 1 -786
box 0 0 112 758
use nand2  g627
timestamp 1543772396
transform 1 0 5768 0 1 -786
box 0 0 112 758
use nand2  g617
timestamp 1543772396
transform 1 0 5880 0 1 -786
box 0 0 112 758
use nand2  g622
timestamp 1543772396
transform 1 0 5992 0 1 -786
box 0 0 112 758
use nand2  g613
timestamp 1543772396
transform 1 0 6104 0 1 -786
box 0 0 112 758
use nand2  g612
timestamp 1543772396
transform 1 0 6216 0 1 -786
box 0 0 112 758
use nand2  g611
timestamp 1543772396
transform 1 0 6328 0 1 -786
box 0 0 112 758
use nand2  g616
timestamp 1543772396
transform 1 0 6440 0 1 -786
box 0 0 112 758
use nand2  g625
timestamp 1543772396
transform 1 0 6552 0 1 -786
box 0 0 112 758
use nand2  g628
timestamp 1543772396
transform 1 0 6664 0 1 -786
box 0 0 112 758
use nand2  g623
timestamp 1543772396
transform 1 0 6776 0 1 -786
box 0 0 112 758
use inv  g630
timestamp 1543772090
transform 1 0 6888 0 1 -786
box 0 0 84 758
use inv  g624
timestamp 1543772090
transform 1 0 6972 0 1 -786
box 0 0 84 758
use inv  g635
timestamp 1543772090
transform 1 0 7056 0 1 -786
box 0 0 84 758
use inv  g631
timestamp 1543772090
transform 1 0 7140 0 1 -786
box 0 0 84 758
use inv  g636
timestamp 1543772090
transform 1 0 7224 0 1 -786
box 0 0 84 758
use nand2  g632
timestamp 1543772396
transform 1 0 7308 0 1 -786
box 0 0 112 758
use nand2  g634
timestamp 1543772396
transform 1 0 7420 0 1 -786
box 0 0 112 758
use nand3  g629
timestamp 1543772418
transform 1 0 7532 0 1 -786
box 0 0 140 758
use nand2  g639
timestamp 1543772396
transform 1 0 7672 0 1 -786
box 0 0 112 758
use nand2  g640
timestamp 1543772396
transform 1 0 7784 0 1 -786
box 0 0 112 758
use nand2  g633
timestamp 1543772396
transform 1 0 7896 0 1 -786
box 0 0 112 758
use nand2  g638
timestamp 1543772396
transform 1 0 8008 0 1 -786
box 0 0 112 758
use nand2  g637
timestamp 1543772396
transform 1 0 8120 0 1 -786
box 0 0 112 758
use inv  g645
timestamp 1543772090
transform 1 0 8232 0 1 -786
box 0 0 84 758
use rightend  rightend_0
timestamp 1544089828
transform 1 0 8316 0 1 -786
box 0 0 308 758
<< labels >>
rlabel metal1 0 28 0 38 3 Done
rlabel metal1 0 56 0 66 3 Req
rlabel metal1 0 84 0 94 3 SDO
rlabel metal2 140 -1388 152 -1388 1 SDI
rlabel metal2 168 -1388 180 -1388 1 Test
rlabel metal2 196 -1388 208 -1388 1 Clock
rlabel metal2 224 -1388 236 -1388 1 nReset
rlabel metal2 252 -1388 264 -1388 1 Load
rlabel metal2 280 -1388 292 -1388 1 nZ
rlabel metal2 308 -1388 320 -1388 1 nBorrow
rlabel metal2 336 -1388 348 -1388 1 LoadAcc
rlabel metal2 364 -1388 376 -1388 1 LoadResult
rlabel metal2 392 -1388 404 -1388 1 ShiftIn
<< end >>
